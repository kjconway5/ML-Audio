module log_lut #(
    parameter int ACCUM_W   = 54,
    parameter int N_MELS    = 40,
    parameter int LOG_OUT_W = 16,
    parameter int LUT_FRAC  = 6,
    parameter int Q_FRAC    = 12
)(
    input  logic                              clk,
    input  logic                              reset,

    // from mel_filterbank
    input  logic [ACCUM_W-1:0]               mel_energy_i [N_MELS],

    // from frame_controller
    input  logic [$clog2(N_MELS)-1:0]        mel_idx_i,
    input  logic                              log_en_i,

    // to output_buffer
    output logic [LOG_OUT_W-1:0]             log_out_o [N_MELS],
    output logic                             log_done_o
);

    // LUT ROM
    // 64 entries, stores log2(1 + frac) in Q4.12
    // generated by python script, ../data/log2_lut.hex
    // TODO: replace with case statement for ASIC synthesis
    logic [LOG_OUT_W-1:0] lut_mem [0:(1<<LUT_FRAC)-1];
    initial $readmemh("../data/log2_lut.hex", lut_mem);

    // select curr mel energy
    logic [ACCUM_W-1:0] current_energy;
    assign current_energy = mel_energy_i[mel_idx_i];

    // PULP IP to compute floor(log2(cur_energy))
    logic [$clog2(ACCUM_W)-1:0] log2_int;

    Log2 #(
        .width(ACCUM_W),
        .speed(2)
    ) u_log2 (
        .A(current_energy),
        .Z(log2_int)
    );

    // Fractional part with LUT
    // extract LUT_FRAC bits just below the leading 1 bit
    // these index into the LUT to get log2(1 + frac)
    logic [LUT_FRAC-1:0]  lut_addr;
    logic [LOG_OUT_W-1:0] lut_val;

    assign lut_addr = (log2_int >= LUT_FRAC)
                    ? current_energy >> (log2_int - LUT_FRAC)
                    : current_energy << (LUT_FRAC - log2_int);

    assign lut_val = lut_mem[lut_addr];

    // Combine integer and fractional parts
    // integer part in Q4.12: floor(log2(x)) shifted left by Q_FRAC
    // fractional part: lut_val already in Q4.12
    // full result = integer + fractional
    logic [LOG_OUT_W-1:0] log_result;

    assign log_result = (current_energy == '0)
                      ? '0
                      : (log2_int << Q_FRAC) + lut_val;

    // Register Output
    // each cycle log_en is high, write result for current mel_idx
    // takes 40 cycles total to compress all mel bins
    // fires log_done_o on the cycle the last bin is written
    always_ff @(posedge clk) begin
        if (reset) begin
            log_done_o <= 1'b0;
            for (int i = 0; i < N_MELS; i++)
                log_out_o[i] <= '0;
        end else begin
            log_done_o <= 1'b0;

            if (log_en_i) begin
                log_out_o[mel_idx_i] <= log_result;

                if (mel_idx_i == N_MELS-1)
                    log_done_o <= 1'b1;
            end
        end
    end

endmodule