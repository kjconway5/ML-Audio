module hpf (#()
    input  logic        clk,
    input  logic        rst_n,
    input  logic [15:0] in_data,
    output logic [15:0] out_data
);


endmodule
