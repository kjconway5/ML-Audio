// Author: Kye Conway

module fir (
    input clk,
    input rst,
    

);



endmodule