module stfft #(
    parameter IW = 16,
    parameter OW = 18,
    parameter FFT_SIZE = 256,
    parameter HOP_SIZE = 128 
)(
    input  wire             i_clk,
    input  wire             i_reset,
    input  wire             i_ce,
    input  wire [IW-1:0]    i_sample,
    output wire [2*OW-1:0]  o_fft_result,
    output wire             o_fft_sync
);

    // Add i_alt_ce logic

    wire [IW-1:0]    win_sample,
    // Windowing
    windowfn #(
        .IW(IW),
        .OW(OW),
        .TW(IW),
        .LGNFFT($clog2(FFT_SIZE))
        /*TODO*/
        /* hanning.hex */
    ) win (
        .i_clk(i_clk),
        .i_reset(i_reset),
        .i_tap_wr(1'b0),
        .i_tap({IW{1'b0}}),
        .i_ce(i_ce),
        .i_alt_ce(/*TODO*/),
        .i_sample(i_sample),
        .o_sample(win_sample),
        .o_ce(win_ce),
        .o_frame()
    );

    // FFT
    fftmain fft (
        .i_clk(i_clk),
        .i_reset(i_reset),
        .i_ce(win_ce),
        .i_sample({win_sample, {IW{1'b0}}}), // real + 0 imaginary
        .o_result(o_fft_result),
        .o_sync(o_fft_sync)
    );



endmodule
